module Top;
//연결 변수 선언
reg[3:0]A,B;
reg C_IN;
wire[3:0] SUM;
wire C_OUT;

endmodule