module fulladd4(output reg[3:0] sum, ouput reg c_out, input [3:0] a,b,input c_in);
//포트 목록만 나열하고 내부에 선언할 수도 있지만 위와 같이 한줄에 포트 선언까지 다 해도 됨
endmodule