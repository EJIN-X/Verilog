//포트는 모듈이 외부 환경과 소통할 수 있는 인터페이스
module fulladd4(sum,c_out,a,b,c_in);
module Top;